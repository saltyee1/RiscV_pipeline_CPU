module Forwarding_Unit(
	input [4:0] D_E_rs1_index,
	input [4:0] D_E_rs2_index,
	input [4:0] E_M_rd_index,
	input [4:0] M_W_rd_index,
	output reg rs1_sel,
	output reg rs2_sel
);
parameter not_forward = 2'd0;
parameter forward_M = 2'd1;
parameter forward_W = 2'd2;
always@(*) begin
	if (D_E_rs1_index == E_M_rd_index)
		rs1_sel = forward_M;
	else if (D_E_rs1_index == M_W_rd_index)
		rs1_sel = forward_W;
	else 
		rs1_sel = not_forward;
end

always@(*) begin
	if (D_E_rs2_index == E_M_rd_index)
		rs2_sel = forward_M;
	else if (D_E_rs2_index == M_W_rd_index)
		rs2_sel = forward_W;
	else 
		rs2_sel = not_forward;
end

endmodule
